dependent source #2  (20110927)

*  + -
V1 1 0 DC 20
R1 1 2 1k

VSENS 66 2 DC 0
R2 66 0 2k

*  - +
F1 3 4 VSENS 3.0 
R3 2 3 3k
R4 3 0 4k
R5 3 4 5k
R6 4 0 6k

* ISC - short circuit current
VSC 4 0 DC 0

.DC V1 20 20 1
*.PRINT DC V(2), V(3), V(4)
.PRINT DC I(VSC)

.END
